import arriskv_pkg::*;

module arriskv_tb;

endmodule